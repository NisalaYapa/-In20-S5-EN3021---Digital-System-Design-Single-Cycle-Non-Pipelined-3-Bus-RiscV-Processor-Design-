module instructionmemory #(parameter Width = 32)(
    input clk,
    input [Width-1:0] address,
	 input MemCopy1,
	 input mul,
    output [Width-1:0] RD
    );
	reg [Width-1:0] mem1[511:0];
	reg MemEn;
	reg [31:0] tempRD;

	initial
	begin
	MemEn = 0;
	tempRD = mem1[0];
	
	
	//mem1[0] = 32'b00000000001000010000001000010011;       	 // ADDI  000000000010 00010 000 00100 0010011
	mem1[0] = 32'b00000000110100011000001010000011;		       //LB     000000001101 00011 000 00101 0000011
	mem1[4] = 32'b00000000001000010000001000010011;       	 // ADDI  000000000011 00010 000 00101 0010011
	
	mem1[8] = 32'b00000000010100100000001010110011;    //add                0000000 00101 00100 000 00101 0110011
   mem1[12] = 32'b01000000010100100000001010110011;   //sub                0100000 00101 00100 000 00101 0110011	
	mem1[16] = 32'b00000000010100100000001010110011;   //add                0000000 00101 00100 000 00101 0110011
	
	
	                            

		// R type                                                                       r1    r2       r3
//		mem1[0] = 32'b00000000001000001000001000110011;   //add                0000000 00010 00001 000 00100 0110011
//		mem1[4] = 32'b01000000001100001000001100110011;   //sub                0100000 00011 00001 000 00110 0110011
//		mem1[8] = 32'b00000000001000001001001010110011;   //SLL                0000000 00010 00001 001 00101 0110011
//		mem1[12] = 32'b00000000001000110010001100110011;  //SLT                0000000 00010 00110 010 00110 0110011
//		mem1[16] = 32'b00000000001100011011000010110011;  //SLTU               0000000 00011 00011 011 00001 0110011
		mem1[20] = 32'b00000000011000011100001010110011;  // XOR               0000000 00110 00011 100 00101 0110011
		mem1[24] = 32'b00000000000100101101001100110011;  // SRL               0000000 00001 00101 101 00110 0110011
		mem1[28] = 32'b01000000011000001101001010110011;  // SRA               0100000 00110 00001 101 00101 0110011
		mem1[32] = 32'b00000000001100001110001110110011;  // OR                0000000 00011 00001 110 00111 0110011
		mem1[36] = 32'b00000000001000011111000010110011;  // AND               0000000 00010 00011 111 00001 0110011

		//I type
																						//      Immediate    R1        Rd
		mem1[40] = 32'b00000000001100010000001000010011;       	// ADDI  000000000011 00010 000 00100 0010011
		mem1[44] = 32'b00000000001100011010001000010011;			// SLTI  000000000011 00011 010 00100 0010011
		mem1[48] = 32'b00000000001100110011001000010011;			//SLTIU  000000000011 00110 011 00100 0010011
		mem1[52] = 32'b00000000001101010100001000010011;			//XORI   000000000011 01010 100 00100 0010011
		mem1[56] = 32'b00000000001100010110001000010011;			//ORI    000000000011 00010 110 00100 0010011
		mem1[60] = 32'b00000000001100110111001000010011;			//ANDI   000000000011 00110 111 00100 0010011
		mem1[64] = 32'b00000000001100011001001000010011;			//SLLI   000000000011 00011 001 00100 0010011
		mem1[68] = 32'b00000000001101000101001000010011;			//SRLI   000000000011 01000 101 00100 0010011
		mem1[72] = 32'b01000000001100010101001000010011;			//SRAI   010000000011 00010 101 00100 0010011


		//S type
																				//      imm1    r2     r1      imm2
		mem1[76] = 32'b00000010001100100000001110100011;		//SB  0000001 00011 00100 000 00111 0100011
		mem1[80] = 32'b00000100001000100001001110100011;		//SH  0000010 00010 00100 001 00111 0100011
		mem1[84] = 32'b00000110011000100010001110100011;		//SW  0000011 00110 00100 010 00111 0100011

		//Sb type

		mem1[88] = 32'b00000110000100001000000011100011;		//BEQ 	 0000011 00001 00001 000 00001 1100011
		mem1[92] = 32'b00000110000100011000000011100011;		//BEQ 	 0000011 00001 00011 000 00001 1100011

		mem1[96] = 32'b00000110000100001001000011100011;		//BNE 	 0000011 00001 00001 001 00001 1100011
		mem1[100] = 32'b00000110000100011001000011100011;		//BNE 	 0000011 00001 00011 001 00001 1100011

		mem1[104] = 32'b00000110000100001100000011100011;		//BLT		 0000011 00001 00001 100 00001 1100011
		mem1[108] = 32'b00000110000100011100000011100011;		//BLT		 0000011 00001 00011 100 00001 1100011

		mem1[112] = 32'b00000110000100001101000011100011;		//BGE		 0000011 00001 00001 101 00001 1100011
		mem1[116] = 32'b00000110000100011101000011100011;		//BGE		 0000011 00001 00011 101 00001 1100011

		mem1[120] = 32'b00000110000100001110000011100011;		//BLTU	 0000011 00001 00001 110 00001 1100011
		mem1[124] = 32'b00000110000100011110000011100011;		//BLTU	 0000011 00001 00011 110 00001 1100011

		mem1[128] = 32'b00000110000100001111000011100011;		//BGEU	 0000011 00001 00001 111 00001 1100011
		mem1[132] = 32'b00000110000100011111000011100011;		//BGEU	 0000011 00001 00011 111 00001 1100011


		//Lw - instuctions
																				//        Imm         r1        rd
		mem1[136] = 32'b00000000110100011000001010000011;		//LB   000000001101 00011 000 00101 0000011
		mem1[140] = 32'b00000000110100111001001010000011;		//LH	 000000001101 00111 001 00101 0000011
		mem1[144] = 32'b00000000110100001010001010000011;		//LW   000000001101 00001 010 00101 0000011
		mem1[148] = 32'b00000000110100010100001010000011;		//LBU  000000001101 00010 100 00101 0000011
		mem1[152] = 32'b00000000110101001101001010000011;		//LHU  000000001101 01001 101 00101 0000011

      /*
		// MEMCOPY
																			  //  Base mem     N        rd   opcode
		mem1[156] = 32'b00000000011100100110000101000000;  // 000000000111 00100 110 00010 1000000
																	//offset 000000000001 00000 000 00001 0000000

		
		mem1[160] = 32'b00000000110100011000001010000011;		//LB   000000001101 00011 000 00101 0000011
		mem1[164] = 32'b00000000110100111001001010000011;		//LH	 000000001101 00111 001 00101 0000011
		mem1[168] = 32'b00000000110100001010001010000011;		//LW   000000001101 00001 010 00101 0000011
		mem1[172] = 32'b00000000110100010100001010000011;		//LBU  000000001101 00010 100 00101 0000011
		mem1[176] = 32'b00000000110101001101001010000011;		//LHU  000000001101 01001 101 00101 0000011

		//MUL                                               //               R1    R2        R3
		mem1[180] = 32'b00000000001000101000001001111111;   // MUL 0000000 00010 00101 000 00100 1111111
		

		mem1[184] = 32'b00000000110100011000001010000011;		//LB   000000001101 00011 000 00101 0000011
		mem1[188] = 32'b00000000110100111001001010000011;		//LH	 000000001101 00111 001 00101 0000011
		mem1[192] = 32'b00000000110100001010001010000011;		//LW   000000001101 00001 010 00101 0000011
		mem1[196] = 32'b00000000110100010100001010000011;		//LBU  000000001101 00010 100 00101 0000011
		mem1[200] = 32'b00000000110101001101001010000011;		//LHU  000000001101 01001 101 00101 0000011
		*/
	end

	always @(MemCopy1) begin
			if(MemCopy1 == 1)
				MemEn = 1;
			if(MemCopy1 == 0)
				MemEn = 0;
		end

	always @(posedge clk) begin
		if(MemEn == 0)
			begin
				tempRD <= mem1[address];     // General instructions
			end
		else
			begin
				if(mul == 1)
					begin
						tempRD <= RD;         // MUL instructions
					end 
				else
					begin
						tempRD <= RD +32'b00000000000100000000000010000000;    // MemCopy instructions
					end
			end
	end
	assign RD = tempRD;


endmodule
